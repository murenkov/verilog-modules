module or_gate(
    input   a,
    input   b,

    output  result
);

assign result = a | b;

endmodule
