module inverse(
    input data,

    output result
);

    assign result = ~data;

endmodule

